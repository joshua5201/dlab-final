`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:36:18 01/07/2016 
// Design Name: 
// Module Name:    GP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module GP(input clk, input reset, input [9:0] x, input [9:0] y, input [9:0] position_x, input [1:0] state, output reg [2:0] rgb);
localparam INIT = 2'd0, GAME = 2'd1, WAIT = 2'd2;
reg [31:0] gp_col;

reg open;
reg [31:0] clk_count;
always @(posedge clk)
begin
	if (reset) begin
		clk_count <= 0;
		open <= 1;
	end
	else begin
		if (clk_count < 5000000) begin
			open <= 1;
			clk_count <= clk_count + 1;
		end
		else if (clk_count >= 5000000 && clk_count <= 10000000) begin
			open <= 0;
			clk_count <= clk_count + 1;
		end
		else if (clk_count > 10000000) begin
			clk_count <= 0;
		end
		else begin
		end
	end
end

always @(*) begin
	if (state == GAME && x - position_x < 32 && x - position_x >= 0 && y > 448) begin
		case (x - position_x)
			0: rgb = gp_col[31] ? 3'b110 : 3'b000;
			1: rgb = gp_col[30] ? 3'b110 : 3'b000;
			2: rgb = gp_col[29] ? 3'b110 : 3'b000;
			3: rgb = gp_col[28] ? 3'b110 : 3'b000;
			4: rgb = gp_col[27] ? 3'b110 : 3'b000;
			5: rgb = gp_col[26] ? 3'b110 : 3'b000;
			6: rgb = gp_col[25] ? 3'b110 : 3'b000;
			7: rgb = gp_col[24] ? 3'b110 : 3'b000;
			8: rgb = gp_col[23] ? 3'b110 : 3'b000;
			9: rgb = gp_col[22] ? 3'b110 : 3'b000;
		 10: rgb = gp_col[21] ? 3'b110 : 3'b000;
		 11: rgb = gp_col[20] ? 3'b110 : 3'b000;
		 12: rgb = gp_col[19] ? 3'b110 : 3'b000;
		 13: rgb = gp_col[18] ? 3'b110 : 3'b000;
		 14: rgb = gp_col[17] ? 3'b110 : 3'b000;
		 15: rgb = gp_col[16] ? 3'b110 : 3'b000;
		 16: rgb = gp_col[15] ? 3'b110 : 3'b000;
		 17: rgb = gp_col[14] ? 3'b110 : 3'b000;
		 18: rgb = gp_col[13] ? 3'b110 : 3'b000;
		 19: rgb = gp_col[12] ? 3'b110 : 3'b000;
		 20: rgb = gp_col[11] ? 3'b110 : 3'b000;
		 21: rgb = gp_col[10] ? 3'b110 : 3'b000;
		 22: rgb = gp_col[9] ? 3'b110 : 3'b000;
		 23: rgb = gp_col[8] ? 3'b110 : 3'b000;
		 24: rgb = gp_col[7] ? 3'b110 : 3'b000;
		 25: rgb = gp_col[6] ? 3'b110 : 3'b000;
		 26: rgb = gp_col[5] ? 3'b110 : 3'b000;
		 27: rgb = gp_col[4] ? 3'b110 : 3'b000;
		 28: rgb = gp_col[3] ? 3'b110 : 3'b000;
		 29: rgb = gp_col[2] ? 3'b110 : 3'b000;
		 30: rgb = gp_col[1] ? 3'b110 : 3'b000;
		 31: rgb = gp_col[0] ? 3'b110 : 3'b000;
		 default: rgb = 3'b000;
		endcase
	end
	else begin
		rgb = 3'b000;
	end
end

always @(*) begin
	if (open) begin
	case (y - 448) 
		 0: gp_col = 32'b00000000000000000000000000000000;
		 1: gp_col = 32'b00000000000000000000000000000000;
		 2: gp_col = 32'b00000000000000000000000000000000;
		 3: gp_col = 32'b00011000000000000000000000001000;
		 4: gp_col = 32'b00011100000000000000000000011000;
		 5: gp_col = 32'b00111111000000000000000011111100;
		 6: gp_col = 32'b00111111000000000000000011111100;
		 7: gp_col = 32'b00111111100000000000000011111100;
		 8: gp_col = 32'b00111111110000000000001111111100;
		 9: gp_col = 32'b01111111111000000000001111111110;
	  10: gp_col = 32'b01111111111100000000011111111110;
		11: gp_col = 32'b01111111111110000000111111111110;
		12: gp_col = 32'b01111111111111000001111111111110;
		13: gp_col = 32'b01111111111111100011111111111110;
		14: gp_col = 32'b11111111111111110111111111111111;
		15: gp_col = 32'b11111111111111111111111111111111;
		16: gp_col = 32'b11111111111111111111111111111111;
		17: gp_col = 32'b01111111111111111111111111111110;
		18: gp_col = 32'b01111111111111111111111111111110;
		19: gp_col = 32'b01111111111111111111111111111110;
		20: gp_col = 32'b01111111111111111111111111111110;
		21: gp_col = 32'b01111111111111111111111111111110;
		22: gp_col = 32'b00111111111111111111111111111100;
		23: gp_col = 32'b00111111111111111111111111111100;
		24: gp_col = 32'b00111111111111111111111111111100;
		25: gp_col = 32'b00111111111111111111111111111100;
		26: gp_col = 32'b00011111111111111111111111111000;
		27: gp_col = 32'b00001111111111111111111111110000;
		28: gp_col = 32'b00000111111111111111111111100000;
		29: gp_col = 32'b00000011111111111111111111000000;
		30: gp_col = 32'b00000001111111111111111110000000;
		31: gp_col = 32'b00000000000011111111000000000000;
		default: gp_col = 32'd0;
	endcase
	end
	else begin
	case (y - 448) 
		 0: gp_col = 32'b00000000000111111111110000000000;
		 1: gp_col = 32'b00000011111111111111111111000000;
		 2: gp_col = 32'b00000111111111111111111111000000;
		 3: gp_col = 32'b00011111111111111111111111111000;
		 4: gp_col = 32'b00011111111111111111111111111000;
		 5: gp_col = 32'b00111111111111111111111111111100;
		 6: gp_col = 32'b00111111111111111111111111111100;
		 7: gp_col = 32'b00111111111111111111111111111100;
		 8: gp_col = 32'b00111111111111111111111111111100;
		 9: gp_col = 32'b01111111111111111111111111111110;
	  10: gp_col = 32'b01111111111111111111111111111110;
		11: gp_col = 32'b01111111111111111111111111111110;
		12: gp_col = 32'b01111111111111111111111111111110;
		13: gp_col = 32'b01111111111111111111111111111110;
		14: gp_col = 32'b11111111111111111111111111111111;
		15: gp_col = 32'b11111111111111111111111111111111;
		16: gp_col = 32'b11111111111111111111111111111111;
		17: gp_col = 32'b01111111111111111111111111111110;
		18: gp_col = 32'b01111111111111111111111111111110;
		19: gp_col = 32'b01111111111111111111111111111110;
		20: gp_col = 32'b01111111111111111111111111111110;
		21: gp_col = 32'b01111111111111111111111111111110;
		22: gp_col = 32'b00111111111111111111111111111100;
		23: gp_col = 32'b00111111111111111111111111111100;
		24: gp_col = 32'b00111111111111111111111111111100;
		25: gp_col = 32'b00111111111111111111111111111100;
		26: gp_col = 32'b00011111111111111111111111111000;
		27: gp_col = 32'b00001111111111111111111111110000;
		28: gp_col = 32'b00000111111111111111111111100000;
		29: gp_col = 32'b00000011111111111111111111000000;
		30: gp_col = 32'b00000001111111111111111110000000;
		31: gp_col = 32'b00000000000011111111000000000000;
		default: gp_col = 32'd0;
	endcase
	end
end

endmodule
